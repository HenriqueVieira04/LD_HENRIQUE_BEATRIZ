-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
-- CREATED		"Thu Sep 19 14:16:21 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY display7 IS 
	PORT
	(
		SW3 :  IN  STD_LOGIC;
		SW2 :  IN  STD_LOGIC;
		SW1 :  IN  STD_LOGIC;
		SW0 :  IN  STD_LOGIC;
		as :  OUT  STD_LOGIC;
		cs :  OUT  STD_LOGIC;
		es :  OUT  STD_LOGIC;
		gs :  OUT  STD_LOGIC;
		fs :  OUT  STD_LOGIC;
		ds :  OUT  STD_LOGIC;
		bs :  OUT  STD_LOGIC
	);
END display7;

ARCHITECTURE bdf_type OF display7 IS 

SIGNAL	A :  STD_LOGIC;
SIGNAL	AN :  STD_LOGIC;
SIGNAL	B :  STD_LOGIC;
SIGNAL	BN :  STD_LOGIC;
SIGNAL	C :  STD_LOGIC;
SIGNAL	CN :  STD_LOGIC;
SIGNAL	D :  STD_LOGIC;
SIGNAL	DN :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_6 <= AN AND BN AND C AND DN;


SYNTHESIZED_WIRE_17 <= AN AND BN AND C;


SYNTHESIZED_WIRE_18 <= AN AND B AND C AND D;


SYNTHESIZED_WIRE_20 <= A AND B AND CN AND DN;


SYNTHESIZED_WIRE_19 <= AN AND BN AND CN;


SYNTHESIZED_WIRE_4 <= A AND B AND DN;


SYNTHESIZED_WIRE_5 <= A AND B AND C;


SYNTHESIZED_WIRE_9 <= B AND C AND D;


SYNTHESIZED_WIRE_12 <= BN AND CN AND D;


SYNTHESIZED_WIRE_13 <= AN AND B AND CN;


SYNTHESIZED_WIRE_11 <= AN AND D;


SYNTHESIZED_WIRE_16 <= AN AND C AND D;


SYNTHESIZED_WIRE_15 <= AN AND BN AND D;


SYNTHESIZED_WIRE_21 <= AN AND B AND CN AND DN;


SYNTHESIZED_WIRE_24 <= AN AND BN AND CN AND D;


SYNTHESIZED_WIRE_22 <= A AND B AND CN AND D;


SYNTHESIZED_WIRE_23 <= A AND BN AND C AND D;


bs <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2 OR SYNTHESIZED_WIRE_3;


SYNTHESIZED_WIRE_0 <= AN AND B AND CN AND D;


SYNTHESIZED_WIRE_3 <= A AND B AND DN;


SYNTHESIZED_WIRE_1 <= B AND C AND DN;


SYNTHESIZED_WIRE_2 <= A AND C AND D;


cs <= SYNTHESIZED_WIRE_4 OR SYNTHESIZED_WIRE_5 OR SYNTHESIZED_WIRE_6;


ds <= SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_7 <= AN AND B AND CN AND DN;


SYNTHESIZED_WIRE_10 <= AN AND BN AND CN AND D;


SYNTHESIZED_WIRE_8 <= A AND BN AND C AND DN;


es <= SYNTHESIZED_WIRE_11 OR SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13;


fs <= SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_15 OR SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_17;


SYNTHESIZED_WIRE_14 <= A AND B AND CN AND D;


gs <= SYNTHESIZED_WIRE_18 OR SYNTHESIZED_WIRE_19 OR SYNTHESIZED_WIRE_20;


AN <= NOT(A);



BN <= NOT(B);



CN <= NOT(C);



DN <= NOT(D);



as <= SYNTHESIZED_WIRE_21 OR SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23 OR SYNTHESIZED_WIRE_24;

A <= SW3;
B <= SW2;
C <= SW1;
D <= SW0;

END bdf_type;